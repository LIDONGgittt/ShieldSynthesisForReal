module design(clock,
  hready, hbusreq0, hlock0, hbusreq1, hlock1, hburst0, hburst1,
  hmaster0, hmastlock, start, decide, locked, hgrant0, hgrant1, busreq, stateA1, stateG2, stateG2_0, stateG2_1, stateG3_0, stateG3_1, stateG3_2, stateG10_1, jx_0, jx_1);

  input clock;
  input hready;
  input hbusreq0;
  input hlock0;
  input hbusreq1;
  input hlock1;
  input hburst0;
  input hburst1;
  output hmaster0;
  output hmastlock;
  output start;
  output decide;
  output locked;
  output hgrant0;
  output hgrant1;
  output busreq;
  output stateA1;
  output stateG2;
  output stateG2_0;
  output stateG2_1;
  output stateG3_0;
  output stateG3_1;
  output stateG3_2;
  output stateG10_1;
  output jx_0;
  output jx_1;
  wire zero;
  wire one;
  wire tmp0;
  wire tmp1;
  wire tmp2;
  wire tmp3;
  wire tmp4;
  wire tmp5;
  wire tmp6;
  wire tmp7;
  wire tmp8;
  wire tmp9;
  wire tmp10;
  wire tmp11;
  wire tmp12;
  wire tmp13;
  wire tmp14;
  wire tmp15;
  wire tmp16;
  wire tmp17;
  wire tmp18;
  wire tmp19;
  wire tmp20;
  wire tmp21;
  wire tmp22;
  wire tmp23;
  wire tmp24;
  wire tmp25;
  wire tmp26;
  wire tmp27;
  wire tmp28;
  wire tmp29;
  wire tmp30;
  wire tmp31;
  wire tmp32;
  wire tmp33;
  wire tmp34;
  wire tmp35;
  wire tmp36;
  wire tmp37;
  wire tmp38;
  wire tmp39;
  wire tmp40;
  wire tmp41;
  wire tmp42;
  wire tmp43;
  wire tmp44;
  wire tmp45;
  wire tmp46;
  wire tmp47;
  wire tmp48;
  wire tmp49;
  wire tmp50;
  wire tmp51;
  wire tmp52;
  wire tmp53;
  wire tmp54;
  wire tmp55;
  wire tmp56;
  wire tmp57;
  wire tmp58;
  wire tmp59;
  wire tmp60;
  wire tmp61;
  wire tmp62;
  wire tmp63;
  wire tmp64;
  wire tmp65;
  wire tmp66;
  wire tmp67;
  wire tmp68;
  wire tmp69;
  wire tmp70;
  wire tmp71;
  wire tmp72;
  wire tmp73;
  wire tmp74;
  wire tmp75;
  wire tmp76;
  wire tmp77;
  wire tmp78;
  wire tmp79;
  wire tmp80;
  wire tmp81;
  wire tmp82;
  wire tmp83;
  wire tmp84;
  wire tmp85;
  wire tmp86;
  wire tmp87;
  wire tmp88;
  wire tmp89;
  wire tmp90;
  wire tmp91;
  wire tmp92;
  wire tmp93;
  wire tmp94;
  wire tmp95;
  wire tmp96;
  wire tmp97;
  wire tmp98;
  wire tmp99;
  wire tmp100;
  wire tmp101;
  wire tmp102;
  wire tmp103;
  wire tmp104;
  wire tmp105;
  wire tmp106;
  wire tmp107;
  wire tmp108;
  wire tmp109;
  wire tmp110;
  wire tmp111;
  wire tmp112;
  wire tmp113;
  wire tmp114;
  wire tmp115;
  wire tmp116;
  wire tmp117;
  wire tmp118;
  wire tmp119;
  wire tmp120;
  wire tmp121;
  wire tmp122;
  wire tmp123;
  wire tmp124;
  wire tmp125;
  wire tmp126;
  wire tmp127;
  wire tmp128;
  wire tmp129;
  wire tmp130;
  wire tmp131;
  wire tmp132;
  wire tmp133;
  wire tmp134;
  wire tmp135;
  wire tmp136;
  wire tmp137;
  wire tmp138;
  wire tmp139;
  wire tmp140;
  wire tmp141;
  wire tmp142;
  wire tmp143;
  wire tmp144;
  wire tmp145;
  wire tmp146;
  wire tmp147;
  wire tmp148;
  wire tmp149;
  wire tmp150;
  wire tmp151;
  wire tmp152;
  wire tmp153;
  wire tmp154;
  wire tmp155;
  wire tmp156;
  wire tmp157;
  wire tmp158;
  wire tmp159;
  wire tmp160;
  wire tmp161;
  wire tmp162;
  wire tmp163;
  wire tmp164;
  wire tmp165;
  wire tmp166;
  wire tmp167;
  wire tmp168;
  wire tmp169;
  wire tmp170;
  wire tmp171;
  wire tmp172;
  wire tmp173;
  wire tmp174;
  wire tmp175;
  wire tmp176;
  wire tmp177;
  wire tmp178;
  wire tmp179;
  wire tmp180;
  wire tmp181;
  wire tmp182;
  wire tmp183;
  wire tmp184;
  wire tmp185;
  wire tmp186;
  wire tmp187;
  wire tmp188;
  wire tmp189;
  wire tmp190;
  wire tmp191;
  wire tmp192;
  wire tmp193;
  wire tmp194;
  wire tmp195;
  wire tmp196;
  wire tmp197;
  wire tmp198;
  wire tmp199;
  wire tmp200;
  wire tmp201;
  wire tmp202;
  wire tmp203;
  wire tmp204;
  wire tmp205;
  wire tmp206;
  wire tmp207;
  wire tmp208;
  wire tmp209;
  wire tmp210;
  wire tmp211;
  wire tmp212;
  wire tmp213;
  wire tmp214;
  wire tmp215;
  wire tmp216;
  wire tmp217;
  wire tmp218;
  wire tmp219;
  wire tmp220;
  wire tmp221;
  wire tmp222;
  wire tmp223;
  wire tmp224;
  wire tmp225;
  wire tmp226;
  wire tmp227;
  wire tmp228;
  wire tmp229;
  wire tmp230;
  wire tmp231;
  wire tmp232;
  wire tmp233;
  wire tmp234;
  wire tmp235;
  wire tmp236;
  wire tmp237;
  wire tmp238;
  wire tmp239;
  wire tmp240;
  wire tmp241;
  wire tmp242;
  wire tmp243;
  wire tmp244;
  wire tmp245;
  wire tmp246;
  wire tmp247;
  wire tmp248;
  wire tmp249;
  wire tmp250;
  wire tmp251;
  wire tmp252;
  wire tmp253;
  wire tmp254;
  wire tmp255;
  wire tmp256;
  wire tmp257;
  wire tmp258;
  wire tmp259;
  wire tmp260;
  wire tmp261;
  wire tmp262;
  wire tmp263;
  wire tmp264;
  wire tmp265;
  wire tmp266;
  wire tmp267;
  wire tmp268;
  wire tmp269;
  wire tmp270;
  wire tmp271;
  wire tmp272;
  wire tmp273;
  wire tmp274;
  wire tmp275;
  wire tmp276;
  wire tmp277;
  wire tmp278;
  wire tmp279;
  wire tmp280;
  wire tmp281;
  wire tmp282;
  wire tmp283;
  wire tmp284;
  wire tmp285;
  wire tmp286;
  wire tmp287;
  wire tmp288;
  wire tmp289;
  wire tmp290;
  wire tmp291;
  wire tmp292;
  wire tmp293;
  wire tmp294;
  wire tmp295;
  wire tmp296;
  wire tmp297;
  wire tmp298;
  wire tmp299;
  wire tmp300;
  wire tmp301;
  wire tmp302;
  wire tmp303;
  wire tmp304;
  wire tmp305;
  wire tmp306;
  wire tmp307;
  wire tmp308;
  wire tmp309;
  wire tmp310;
  wire tmp311;
  wire tmp312;
  wire tmp313;
  wire tmp314;
  wire tmp315;
  wire tmp316;
  wire tmp317;
  wire tmp318;
  wire tmp319;
  wire tmp320;
  wire tmp321;
  wire tmp322;
  wire tmp323;
  wire tmp324;
  wire tmp325;
  wire tmp326;
  wire tmp327;
  wire tmp328;
  wire tmp329;
  wire tmp330;
  wire tmp331;
  wire tmp332;
  wire tmp333;
  wire tmp334;
  wire tmp335;
  wire tmp336;
  wire tmp337;
  wire tmp338;
  wire tmp339;
  wire tmp340;
  wire tmp341;
  wire tmp342;
  wire tmp343;
  wire tmp344;
  wire tmp345;
  wire tmp346;
  wire tmp347;
  wire tmp348;
  wire tmp349;
  wire tmp350;
  wire tmp351;
  wire tmp352;
  wire tmp353;
  wire tmp354;
  wire tmp355;
  wire tmp356;
  wire tmp357;
  wire tmp358;
  wire tmp359;
  wire tmp360;
  wire tmp361;
  wire tmp362;
  wire tmp363;
  wire tmp364;
  wire tmp365;
  wire tmp366;
  wire tmp367;
  wire tmp368;
  wire tmp369;
  wire tmp370;
  wire tmp371;
  wire tmp372;
  wire tmp373;
  wire tmp374;
  wire tmp375;
  wire tmp376;
  wire tmp377;
  wire tmp378;
  wire tmp379;
  wire tmp380;
  wire tmp381;
  wire tmp382;
  wire tmp383;
  wire tmp384;
  wire tmp385;
  wire tmp386;
  wire tmp387;
  wire tmp388;
  wire tmp389;
  wire tmp390;
  wire tmp391;
  wire tmp392;
  wire tmp393;
  wire tmp394;
  wire tmp395;
  wire tmp396;
  wire tmp397;
  wire tmp398;
  wire tmp399;
  wire tmp400;
  wire tmp401;
  wire tmp402;
  wire tmp403;
  wire tmp404;
  wire tmp405;
  wire tmp406;
  wire tmp407;
  wire tmp408;
  wire tmp409;
  wire tmp410;
  wire tmp411;
  wire tmp412;
  wire tmp413;
  wire tmp414;
  wire tmp415;
  wire tmp416;
  wire tmp417;
  wire tmp418;
  wire tmp419;
  wire tmp420;
  wire tmp421;
  wire tmp422;
  wire tmp423;
  wire tmp424;
  wire tmp425;
  wire tmp426;
  wire tmp427;
  wire tmp428;
  wire tmp429;
  wire tmp430;
  wire tmp431;
  wire tmp432;
  wire tmp433;
  wire tmp434;
  wire tmp435;
  wire tmp436;
  wire tmp437;
  wire tmp438;
  wire tmp439;
  wire tmp440;
  wire tmp441;
  wire tmp442;
  wire tmp443;
  wire tmp444;
  wire tmp445;
  wire tmp446;
  wire tmp447;
  wire tmp448;
  wire tmp449;
  wire tmp450;
  wire tmp451;
  wire tmp452;
  wire tmp453;
  wire tmp454;
  wire tmp455;
  wire tmp456;
  wire tmp457;
  wire tmp458;
  wire tmp459;
  wire tmp460;
  wire tmp461;
  wire tmp462;
  wire tmp463;
  wire tmp464;
  wire tmp465;
  wire tmp466;
  wire tmp467;
  wire tmp468;
  wire tmp469;
  wire tmp470;
  wire tmp471;
  wire tmp472;
  wire tmp473;
  wire tmp474;
  wire tmp475;
  wire tmp476;
  wire tmp477;
  wire tmp478;
  wire tmp479;
  wire tmp480;
  wire tmp481;
  wire tmp482;
  wire tmp483;
  wire tmp484;
  wire tmp485;
  wire tmp486;
  wire tmp487;
  wire tmp488;
  wire tmp489;
  wire tmp490;
  wire tmp491;
  wire tmp492;
  wire tmp493;
  wire tmp494;
  wire tmp495;
  wire tmp496;
  wire tmp497;
  wire tmp498;
  wire tmp499;
  wire tmp500;
  wire tmp501;
  wire tmp502;
  wire tmp503;
  wire tmp504;
  wire tmp505;
  wire tmp506;
  wire tmp507;
  wire tmp508;
  wire tmp509;
  wire tmp510;
  wire tmp511;
  wire tmp512;
  wire tmp513;
  wire tmp514;
  wire tmp515;
  wire tmp516;
  wire tmp517;
  wire tmp518;
  wire tmp519;
  wire tmp520;
  wire tmp521;
  wire tmp522;
  wire tmp523;
  wire tmp524;
  wire tmp525;
  wire tmp526;
  wire tmp527;
  wire tmp528;
  wire tmp529;
  wire tmp530;
  wire tmp531;
  wire tmp532;
  wire tmp533;
  wire tmp534;
  wire tmp535;
  wire tmp536;
  wire tmp537;
  wire tmp538;
  wire tmp539;
  wire tmp540;
  wire tmp541;
  wire tmp542;
  wire tmp543;
  wire tmp544;
  wire tmp545;
  wire tmp546;
  wire tmp547;
  wire tmp548;
  wire tmp549;
  wire tmp550;
  wire tmp551;
  wire tmp552;
  wire tmp553;
  wire tmp554;
  wire tmp555;
  wire tmp556;
  wire tmp557;
  wire tmp558;
  wire tmp559;
  wire tmp560;
  wire tmp561;
  wire tmp562;
  wire tmp563;
  wire tmp564;
  wire tmp565;
  wire tmp566;
  wire tmp567;
  wire tmp568;
  wire tmp569;
  wire tmp570;
  wire tmp571;
  wire tmp572;
  wire tmp573;
  wire tmp574;
  wire tmp575;
  wire tmp576;
  wire tmp577;
  wire tmp578;
  wire tmp579;
  wire tmp580;
  wire tmp581;
  wire tmp582;
  wire tmp583;
  wire tmp584;
  wire tmp585;
  wire tmp586;
  wire tmp587;
  wire tmp588;
  wire tmp589;
  wire tmp590;
  wire tmp591;
  wire tmp592;
  wire tmp593;
  wire tmp594;
  wire tmp595;
  wire tmp596;
  wire tmp597;
  wire tmp598;
  wire tmp599;
  wire tmp600;
  wire tmp601;
  wire tmp602;
  wire tmp603;
  wire tmp604;
  wire tmp605;
  wire tmp606;
  wire tmp607;
  wire tmp608;
  wire tmp609;
  wire tmp610;
  wire tmp611;
  wire tmp612;
  wire tmp613;
  wire tmp614;
  wire tmp615;
  wire tmp616;
  wire tmp617;
  wire tmp618;
  wire tmp619;
  wire tmp620;
  wire tmp621;
  wire tmp622;
  wire tmp623;
  wire tmp624;
  wire tmp625;
  wire tmp626;
  wire tmp627;
  wire tmp628;
  wire tmp629;
  wire tmp630;
  wire tmp631;
  wire tmp632;
  wire tmp633;
  wire tmp634;
  wire tmp635;
  wire tmp636;
  wire tmp637;
  wire tmp638;
  wire tmp639;
  wire tmp640;
  wire tmp641;
  wire tmp642;
  wire tmp643;
  wire tmp644;
  wire tmp645;
  wire tmp646;
  wire tmp647;
  wire tmp648;
  wire tmp649;
  wire tmp650;
  wire tmp651;
  wire tmp652;
  wire tmp653;
  wire tmp654;
  wire tmp655;
  wire tmp656;
  wire tmp657;
  wire tmp658;
  wire tmp659;
  wire tmp660;
  wire tmp661;
  wire tmp662;
  wire tmp663;
  wire tmp664;
  wire tmp665;
  wire tmp666;
  wire tmp667;
  wire tmp668;
  wire tmp669;
  wire tmp670;
  wire tmp671;
  wire tmp672;
  wire tmp673;
  wire tmp674;
  wire tmp675;
  wire tmp676;
  wire tmp677;
  wire tmp678;
  wire tmp679;
  wire tmp680;
  wire tmp681;
  wire tmp682;
  wire tmp683;
  wire tmp684;
  wire tmp685;
  wire tmp686;
  wire tmp687;
  wire tmp688;
  wire tmp689;
  wire tmp690;
  wire tmp691;
  wire tmp692;
  wire tmp693;
  wire tmp694;
  wire tmp695;
  wire tmp696;
  wire tmp697;
  wire tmp698;
  wire tmp699;
  wire tmp700;
  wire tmp701;
  wire tmp702;
  wire tmp703;
  wire tmp704;
  wire tmp705;
  wire tmp706;
  wire tmp707;
  wire tmp708;
  wire tmp709;
  wire tmp710;
  wire tmp711;
  wire tmp712;
  wire tmp713;
  wire tmp714;
  wire tmp715;
  wire tmp716;
  wire tmp717;
  wire tmp718;
  wire tmp719;
  wire tmp720;
  wire tmp721;
  wire tmp722;
  wire tmp723;
  wire tmp724;
  wire tmp725;
  wire tmp726;
  wire tmp727;
  wire tmp728;
  wire tmp729;
  wire tmp730;
  wire tmp731;
  wire tmp732;
  wire tmp733;
  wire tmp734;
  wire tmp735;
  wire tmp736;
  wire tmp737;
  wire tmp738;
  wire tmp739;
  wire tmp740;
  wire tmp741;
  wire tmp742;
  wire tmp743;
  wire tmp744;
  wire tmp745;
  wire tmp746;
  wire tmp747;
  wire tmp748;
  wire tmp749;
  wire tmp750;
  wire tmp751;
  wire tmp752;
  wire tmp753;
  wire tmp754;
  wire tmp755;
  wire tmp756;
  wire tmp757;
  wire tmp758;
  wire tmp759;
  wire tmp760;
  wire tmp761;
  wire tmp762;
  wire tmp763;
  wire tmp764;
  wire tmp765;
  wire tmp766;
  wire tmp767;
  wire tmp768;
  wire tmp769;
  wire tmp770;
  wire tmp771;
  wire tmp772;
  wire tmp773;
  wire tmp774;
  wire tmp775;
  wire tmp776;
  wire tmp777;
  wire tmp778;
  wire tmp779;
  wire tmp780;
  wire tmp781;
  wire tmp782;
  wire tmp783;
  wire tmp784;
  wire tmp785;
  wire tmp786;
  wire tmp787;
  wire tmp788;
  wire tmp789;
  reg hready_ps;
  reg hbusreq0_ps;
  reg hlock0_ps;
  reg hbusreq1_ps;
  reg hlock1_ps;
  reg hburst0_ps;
  reg hburst1_ps;
  reg hmaster0_ps;
  reg hmastlock_ps;
  reg start_ps;
  reg decide_ps;
  reg locked_ps;
  reg hgrant0_ps;
  reg hgrant1_ps;
  reg busreq_ps;
  reg stateA1_ps;
  reg stateG2_ps;
  reg stateG2_0_ps;
  reg stateG2_1_ps;
  reg stateG3_0_ps;
  reg stateG3_1_ps;
  reg stateG3_2_ps;
  reg stateG10_1_ps;
  reg jx_0_ps;
  reg jx_1_ps;


  assign tmp0 = hmastlock_ps ? one : zero;
  assign tmp1 = ~tmp0;
  assign tmp2 = start_ps ? one : tmp1;
  assign tmp3 = stateG3_0_ps ? tmp2 : one;
  assign tmp4 = stateG3_1_ps ? tmp3 : one;
  assign tmp5 = stateG3_2_ps ? one : tmp4;
  assign tmp6 = stateG2_ps ? one : tmp5;
  assign tmp7 = stateG3_2_ps ? one : tmp3;
  assign tmp8 = jx_1_ps ? tmp6 : tmp7;
  assign tmp9 = jx_0_ps ? tmp6 : tmp8;
  assign tmp10 = hbusreq1_ps ? tmp6 : tmp9;
  assign tmp11 = hmaster0_ps ? tmp10 : one;
  assign tmp12 = hlock0_ps ? tmp6 : tmp7;
  assign tmp13 = jx_1_ps ? tmp6 : tmp12;
  assign tmp14 = jx_0_ps ? tmp6 : tmp13;
  assign tmp15 = hmaster0_ps ? one : tmp14;
  assign tmp16 = hgrant1_ps ? tmp11 : tmp15;
  assign tmp17 = stateG3_2_ps ? tmp2 : one;
  assign tmp18 = stateG2_ps ? one : tmp17;
  assign tmp19 = jx_1_ps ? tmp18 : tmp17;
  assign tmp20 = jx_0_ps ? tmp18 : tmp19;
  assign tmp21 = hbusreq1_ps ? tmp18 : tmp20;
  assign tmp22 = hbusreq0_ps ? tmp18 : tmp17;
  assign tmp23 = jx_1_ps ? tmp18 : tmp22;
  assign tmp24 = jx_0_ps ? tmp18 : tmp23;
  assign tmp25 = hmaster0_ps ? tmp21 : tmp24;
  assign tmp26 = hlock0_ps ? one : tmp18;
  assign tmp27 = hbusreq0_ps ? tmp26 : tmp18;
  assign tmp28 = hlock0_ps ? one : tmp17;
  assign tmp29 = hbusreq0_ps ? tmp28 : tmp17;
  assign tmp30 = jx_1_ps ? tmp27 : tmp29;
  assign tmp31 = jx_0_ps ? tmp27 : tmp30;
  assign tmp32 = hbusreq1_ps ? tmp18 : tmp31;
  assign tmp33 = hmaster0_ps ? tmp32 : tmp24;
  assign tmp34 = hgrant1_ps ? tmp25 : tmp33;
  assign tmp35 = hready_ps ? tmp16 : tmp34;
  assign tmp36 = stateA1_ps ? tmp6 : tmp5;
  assign tmp37 = busreq_ps ? tmp36 : tmp5;
  assign tmp38 = jx_1_ps ? tmp6 : tmp37;
  assign tmp39 = jx_0_ps ? tmp6 : tmp38;
  assign tmp40 = hmaster0_ps ? tmp39 : one;
  assign tmp41 = hmaster0_ps ? one : tmp39;
  assign tmp42 = hgrant1_ps ? tmp40 : tmp41;
  assign tmp43 = stateA1_ps ? tmp18 : tmp17;
  assign tmp44 = busreq_ps ? tmp43 : tmp17;
  assign tmp45 = jx_1_ps ? tmp18 : tmp44;
  assign tmp46 = jx_0_ps ? tmp18 : tmp45;
  assign tmp47 = hmaster0_ps ? tmp20 : tmp46;
  assign tmp48 = hgrant1_ps ? tmp46 : tmp47;
  assign tmp49 = hready_ps ? tmp42 : tmp48;
  assign tmp50 = decide_ps ? tmp35 : tmp49;
  assign tmp51 = ~tmp50;
  assign tmp52 = hlock1_ps ? one : zero;
  assign tmp53 = locked_ps ? one : zero;
  assign tmp54 = hlock1_ps ? tmp53 : zero;
  assign tmp55 = hlock0_ps ? tmp52 : tmp54;
  assign tmp56 = hburst0_ps ? one : tmp2;
  assign tmp57 = hburst1_ps ? one : tmp56;
  assign tmp58 = ~tmp57;
  assign tmp59 = stateA1_ps ? one : tmp58;
  assign tmp60 = locked_ps ? one : tmp59;
  assign tmp61 = ~tmp60;
  assign tmp62 = hlock1_ps ? one : tmp61;
  assign tmp63 = start_ps ? tmp0 : zero;
  assign tmp64 = stateG3_0_ps ? tmp0 : tmp63;
  assign tmp65 = stateG3_0_ps ? tmp63 : tmp0;
  assign tmp66 = stateG3_1_ps ? tmp64 : tmp65;
  assign tmp67 = stateG3_2_ps ? tmp0 : tmp66;
  assign tmp68 = stateG3_0_ps ? one : tmp2;
  assign tmp69 = stateG3_1_ps ? tmp3 : tmp68;
  assign tmp70 = stateG3_2_ps ? tmp2 : tmp69;
  assign tmp71 = ~tmp70;
  assign tmp72 = hburst0_ps ? tmp67 : tmp71;
  assign tmp73 = ~tmp72;
  assign tmp74 = stateG2_ps ? one : tmp73;
  assign tmp75 = stateA1_ps ? tmp74 : tmp73;
  assign tmp76 = locked_ps ? tmp75 : zero;
  assign tmp77 = hlock1_ps ? tmp76 : zero;
  assign tmp78 = hlock0_ps ? tmp62 : tmp77;
  assign tmp79 = hbusreq0_ps ? tmp78 : tmp54;
  assign tmp80 = hbusreq0_ps ? tmp55 : tmp54;
  assign tmp81 = jx_1_ps ? tmp79 : tmp80;
  assign tmp82 = jx_0_ps ? tmp55 : tmp81;
  assign tmp83 = locked_ps ? one : tmp58;
  assign tmp84 = hlock0_ps ? tmp83 : one;
  assign tmp85 = hbusreq0_ps ? tmp84 : one;
  assign tmp86 = jx_1_ps ? tmp85 : one;
  assign tmp87 = jx_0_ps ? one : tmp86;
  assign tmp88 = ~tmp87;
  assign tmp89 = hbusreq1_ps ? tmp82 : tmp88;
  assign tmp90 = jx_0_ps ? tmp55 : tmp80;
  assign tmp91 = hbusreq1_ps ? tmp90 : zero;
  assign tmp92 = hmaster0_ps ? tmp89 : tmp91;
  assign tmp93 = hlock1_ps ? one : tmp53;
  assign tmp94 = hlock0_ps ? tmp93 : zero;
  assign tmp95 = hbusreq0_ps ? tmp94 : zero;
  assign tmp96 = jx_1_ps ? tmp95 : tmp94;
  assign tmp97 = jx_0_ps ? tmp94 : tmp96;
  assign tmp98 = hlock0_ps ? one : zero;
  assign tmp99 = hbusreq0_ps ? tmp98 : zero;
  assign tmp100 = jx_1_ps ? tmp99 : tmp98;
  assign tmp101 = jx_0_ps ? tmp98 : tmp100;
  assign tmp102 = hbusreq1_ps ? tmp97 : tmp101;
  assign tmp103 = hlock1_ps ? one : tmp76;
  assign tmp104 = hlock1_ps ? tmp60 : one;
  assign tmp105 = ~tmp104;
  assign tmp106 = hlock0_ps ? tmp103 : tmp105;
  assign tmp107 = jx_1_ps ? tmp106 : tmp94;
  assign tmp108 = jx_0_ps ? tmp107 : tmp96;
  assign tmp109 = hbusreq1_ps ? tmp108 : tmp101;
  assign tmp110 = hmaster0_ps ? tmp102 : tmp109;
  assign tmp111 = hgrant1_ps ? tmp92 : tmp110;
  assign tmp112 = hlock1_ps ? tmp0 : zero;
  assign tmp113 = hlock0_ps ? tmp52 : tmp112;
  assign tmp114 = stateA1_ps ? one : tmp0;
  assign tmp115 = ~tmp114;
  assign tmp116 = hlock1_ps ? one : tmp115;
  assign tmp117 = stateG3_1_ps ? tmp2 : tmp3;
  assign tmp118 = stateG3_2_ps ? one : tmp117;
  assign tmp119 = stateG3_1_ps ? tmp0 : tmp64;
  assign tmp120 = stateG3_2_ps ? tmp63 : tmp119;
  assign tmp121 = ~tmp120;
  assign tmp122 = hburst0_ps ? tmp118 : tmp121;
  assign tmp123 = ~tmp122;
  assign tmp124 = stateG2_ps ? tmp0 : tmp123;
  assign tmp125 = stateA1_ps ? tmp124 : tmp123;
  assign tmp126 = hlock1_ps ? tmp125 : zero;
  assign tmp127 = hlock0_ps ? tmp116 : tmp126;
  assign tmp128 = hbusreq0_ps ? tmp127 : tmp112;
  assign tmp129 = hbusreq0_ps ? tmp113 : tmp112;
  assign tmp130 = jx_1_ps ? tmp128 : tmp129;
  assign tmp131 = jx_0_ps ? tmp113 : tmp130;
  assign tmp132 = hlock0_ps ? tmp0 : one;
  assign tmp133 = hbusreq0_ps ? tmp132 : one;
  assign tmp134 = jx_1_ps ? tmp133 : one;
  assign tmp135 = jx_0_ps ? one : tmp134;
  assign tmp136 = ~tmp135;
  assign tmp137 = hbusreq1_ps ? tmp131 : tmp136;
  assign tmp138 = hlock1_ps ? one : tmp125;
  assign tmp139 = busreq_ps ? tmp114 : tmp0;
  assign tmp140 = hlock1_ps ? tmp139 : one;
  assign tmp141 = ~tmp140;
  assign tmp142 = hlock0_ps ? tmp138 : tmp141;
  assign tmp143 = hlock1_ps ? one : tmp0;
  assign tmp144 = hlock0_ps ? tmp143 : zero;
  assign tmp145 = jx_1_ps ? tmp142 : tmp144;
  assign tmp146 = hbusreq0_ps ? tmp144 : zero;
  assign tmp147 = jx_0_ps ? tmp145 : tmp146;
  assign tmp148 = hlock0_ps ? tmp0 : zero;
  assign tmp149 = hbusreq0_ps ? tmp148 : zero;
  assign tmp150 = hbusreq1_ps ? tmp147 : tmp149;
  assign tmp151 = hmaster0_ps ? tmp137 : tmp150;
  assign tmp152 = hbusreq1_ps ? tmp131 : tmp99;
  assign tmp153 = hbusreq1_ps ? tmp147 : tmp99;
  assign tmp154 = hmaster0_ps ? tmp152 : tmp153;
  assign tmp155 = hgrant1_ps ? tmp151 : tmp154;
  assign tmp156 = hready_ps ? tmp111 : tmp155;
  assign tmp157 = decide_ps ? tmp156 : tmp53;
  assign tmp158 = hgrant1_ps ? one : zero;
  assign tmp159 = hmaster0_ps ? one : zero;
  assign tmp160 = hready_ps ? tmp158 : tmp159;
  assign tmp161 = locked_ps ? tmp0 : tmp1;
  assign tmp162 = hmaster0_ps ? tmp161 : zero;
  assign tmp163 = ~tmp161;
  assign tmp164 = hmaster0_ps ? one : tmp163;
  assign tmp165 = ~tmp164;
  assign tmp166 = hgrant1_ps ? tmp162 : tmp165;
  assign tmp167 = hready_ps ? tmp166 : one;
  assign tmp168 = ~tmp167;
  assign tmp169 = hlock1_ps ? tmp53 : one;
  assign tmp170 = hlock0_ps ? one : tmp169;
  assign tmp171 = hburst0_ps ? tmp67 : zero;
  assign tmp172 = hburst1_ps ? tmp72 : tmp171;
  assign tmp173 = hburst0 ? tmp172 : zero;
  assign tmp174 = hburst1 ? tmp172 : tmp173;
  assign tmp175 = ~tmp174;
  assign tmp176 = stateA1_ps ? one : tmp175;
  assign tmp177 = hlock1 ? tmp176 : one;
  assign tmp178 = locked_ps ? tmp177 : zero;
  assign tmp179 = hlock1_ps ? tmp178 : tmp60;
  assign tmp180 = hlock0_ps ? tmp179 : tmp77;
  assign tmp181 = hbusreq0_ps ? tmp180 : tmp53;
  assign tmp182 = hbusreq0_ps ? tmp170 : tmp53;
  assign tmp183 = jx_1_ps ? tmp181 : tmp182;
  assign tmp184 = jx_0_ps ? tmp170 : tmp183;
  assign tmp185 = hbusreq0_ps ? one : zero;
  assign tmp186 = hlock0_ps ? tmp83 : zero;
  assign tmp187 = hbusreq0_ps ? tmp186 : zero;
  assign tmp188 = jx_1_ps ? tmp187 : tmp185;
  assign tmp189 = jx_0_ps ? tmp185 : tmp188;
  assign tmp190 = hbusreq1_ps ? tmp184 : tmp189;
  assign tmp191 = jx_0_ps ? tmp170 : tmp182;
  assign tmp192 = hbusreq1_ps ? tmp191 : tmp185;
  assign tmp193 = hmaster0_ps ? tmp190 : tmp192;
  assign tmp194 = hbusreq0_ps ? tmp93 : one;
  assign tmp195 = jx_1_ps ? tmp194 : tmp93;
  assign tmp196 = jx_0_ps ? tmp93 : tmp195;
  assign tmp197 = hbusreq1_ps ? tmp196 : one;
  assign tmp198 = hlock1_ps ? tmp178 : tmp76;
  assign tmp199 = hlock1_ps ? tmp60 : zero;
  assign tmp200 = hlock0_ps ? tmp198 : tmp199;
  assign tmp201 = jx_1_ps ? tmp200 : tmp93;
  assign tmp202 = jx_0_ps ? tmp201 : tmp195;
  assign tmp203 = hbusreq1_ps ? tmp202 : one;
  assign tmp204 = hmaster0_ps ? tmp197 : tmp203;
  assign tmp205 = ~tmp204;
  assign tmp206 = hgrant1_ps ? tmp193 : tmp205;
  assign tmp207 = hlock1_ps ? tmp0 : one;
  assign tmp208 = hlock0_ps ? one : tmp207;
  assign tmp209 = hburst0_ps ? tmp118 : tmp1;
  assign tmp210 = hburst1_ps ? tmp122 : tmp209;
  assign tmp211 = hburst0 ? tmp210 : tmp1;
  assign tmp212 = hburst1 ? tmp210 : tmp211;
  assign tmp213 = ~tmp212;
  assign tmp214 = stateA1_ps ? tmp0 : tmp213;
  assign tmp215 = hlock1 ? tmp214 : tmp0;
  assign tmp216 = hlock1_ps ? tmp215 : tmp114;
  assign tmp217 = hlock0_ps ? tmp216 : tmp126;
  assign tmp218 = hbusreq0_ps ? tmp217 : tmp0;
  assign tmp219 = hbusreq0_ps ? tmp208 : tmp0;
  assign tmp220 = jx_1_ps ? tmp218 : tmp219;
  assign tmp221 = jx_0_ps ? tmp208 : tmp220;
  assign tmp222 = jx_1_ps ? tmp149 : tmp185;
  assign tmp223 = jx_0_ps ? tmp185 : tmp222;
  assign tmp224 = hbusreq1_ps ? tmp221 : tmp223;
  assign tmp225 = hlock1_ps ? tmp215 : tmp125;
  assign tmp226 = hlock1_ps ? tmp139 : zero;
  assign tmp227 = hlock0_ps ? tmp225 : tmp226;
  assign tmp228 = jx_1_ps ? tmp227 : tmp143;
  assign tmp229 = hbusreq0_ps ? tmp143 : one;
  assign tmp230 = jx_0_ps ? tmp228 : tmp229;
  assign tmp231 = hbusreq0_ps ? tmp0 : one;
  assign tmp232 = hbusreq1_ps ? tmp230 : tmp231;
  assign tmp233 = ~tmp232;
  assign tmp234 = hmaster0_ps ? tmp224 : tmp233;
  assign tmp235 = hbusreq1_ps ? tmp221 : zero;
  assign tmp236 = hbusreq1_ps ? tmp230 : one;
  assign tmp237 = ~tmp236;
  assign tmp238 = hmaster0_ps ? tmp235 : tmp237;
  assign tmp239 = hgrant1_ps ? tmp234 : tmp238;
  assign tmp240 = hready_ps ? tmp206 : tmp239;
  assign tmp241 = decide_ps ? tmp240 : tmp158;
  assign tmp242 = hlock0_ps ? tmp93 : tmp52;
  assign tmp243 = hbusreq0_ps ? tmp242 : one;
  assign tmp244 = jx_1_ps ? tmp243 : tmp242;
  assign tmp245 = jx_0_ps ? tmp242 : tmp244;
  assign tmp246 = hbusreq1_ps ? tmp245 : one;
  assign tmp247 = hmaster0_ps ? tmp246 : tmp203;
  assign tmp248 = ~tmp247;
  assign tmp249 = hgrant1_ps ? tmp193 : tmp248;
  assign tmp250 = hready_ps ? tmp249 : tmp239;
  assign tmp251 = decide_ps ? tmp250 : tmp158;
  assign tmp252 = ~tmp251;
  assign tmp253 = stateG3_2_ps ? tmp2 : tmp117;
  assign tmp254 = stateG2_ps ? one : tmp253;
  assign tmp255 = ~tmp254;
  assign tmp256 = jx_1_ps ? one : tmp255;
  assign tmp257 = jx_1_ps ? one : zero;
  assign tmp258 = ~tmp257;
  assign tmp259 = jx_0_ps ? tmp256 : tmp258;
  assign tmp260 = hlock0_ps ? tmp254 : tmp18;
  assign tmp261 = jx_1_ps ? one : tmp260;
  assign tmp262 = jx_0_ps ? tmp261 : tmp257;
  assign tmp263 = ~tmp260;
  assign tmp264 = jx_1_ps ? one : tmp263;
  assign tmp265 = jx_0_ps ? tmp264 : tmp258;
  assign tmp266 = ~tmp265;
  assign tmp267 = hbusreq1_ps ? tmp262 : tmp266;
  assign tmp268 = ~tmp267;
  assign tmp269 = hmaster0_ps ? tmp259 : tmp268;
  assign tmp270 = ~tmp18;
  assign tmp271 = jx_1_ps ? one : tmp270;
  assign tmp272 = jx_0_ps ? tmp271 : tmp258;
  assign tmp273 = hbusreq1_ps ? tmp259 : tmp272;
  assign tmp274 = jx_1_ps ? one : tmp254;
  assign tmp275 = jx_0_ps ? tmp274 : tmp257;
  assign tmp276 = ~tmp259;
  assign tmp277 = hbusreq1_ps ? tmp275 : tmp276;
  assign tmp278 = ~tmp277;
  assign tmp279 = hmaster0_ps ? tmp273 : tmp278;
  assign tmp280 = hgrant1_ps ? tmp269 : tmp279;
  assign tmp281 = jx_1_ps ? one : tmp18;
  assign tmp282 = jx_0_ps ? tmp281 : tmp257;
  assign tmp283 = ~tmp272;
  assign tmp284 = hbusreq1_ps ? tmp282 : tmp283;
  assign tmp285 = ~tmp284;
  assign tmp286 = hmaster0_ps ? tmp259 : tmp285;
  assign tmp287 = ~tmp17;
  assign tmp288 = jx_1_ps ? one : tmp287;
  assign tmp289 = jx_0_ps ? tmp288 : tmp258;
  assign tmp290 = hbusreq1_ps ? tmp289 : tmp272;
  assign tmp291 = hmaster0_ps ? tmp290 : tmp278;
  assign tmp292 = hgrant1_ps ? tmp286 : tmp291;
  assign tmp293 = decide_ps ? tmp280 : tmp292;
  assign tmp294 = ~tmp293;
  assign tmp295 = ~tmp63;
  assign tmp296 = hburst0_ps ? one : tmp295;
  assign tmp297 = hburst1_ps ? one : tmp296;
  assign tmp298 = ~tmp297;
  assign tmp299 = stateG2_ps ? tmp0 : tmp298;
  assign tmp300 = hbusreq1_ps ? tmp299 : zero;
  assign tmp301 = hmaster0_ps ? tmp300 : zero;
  assign tmp302 = hlock0_ps ? tmp299 : zero;
  assign tmp303 = hbusreq0_ps ? tmp302 : zero;
  assign tmp304 = jx_1_ps ? tmp303 : tmp302;
  assign tmp305 = jx_0_ps ? tmp302 : tmp304;
  assign tmp306 = ~tmp305;
  assign tmp307 = hmaster0_ps ? one : tmp306;
  assign tmp308 = ~tmp307;
  assign tmp309 = hgrant1_ps ? tmp301 : tmp308;
  assign tmp310 = jx_0_ps ? tmp302 : tmp303;
  assign tmp311 = hbusreq1_ps ? tmp310 : tmp303;
  assign tmp312 = hmaster0_ps ? tmp300 : tmp311;
  assign tmp313 = hready_ps ? tmp309 : tmp312;
  assign tmp314 = stateG2_ps ? one : tmp297;
  assign tmp315 = ~tmp314;
  assign tmp316 = busreq_ps ? tmp299 : tmp315;
  assign tmp317 = jx_1_ps ? tmp299 : tmp316;
  assign tmp318 = jx_0_ps ? tmp317 : tmp316;
  assign tmp319 = ~tmp316;
  assign tmp320 = jx_1_ps ? tmp314 : tmp319;
  assign tmp321 = jx_0_ps ? tmp320 : tmp319;
  assign tmp322 = ~tmp321;
  assign tmp323 = hbusreq1_ps ? tmp318 : tmp322;
  assign tmp324 = hmaster0_ps ? tmp323 : zero;
  assign tmp325 = hbusreq0_ps ? tmp299 : tmp315;
  assign tmp326 = jx_1_ps ? tmp325 : tmp316;
  assign tmp327 = jx_0_ps ? tmp316 : tmp326;
  assign tmp328 = ~tmp327;
  assign tmp329 = hmaster0_ps ? one : tmp328;
  assign tmp330 = ~tmp329;
  assign tmp331 = hgrant1_ps ? tmp324 : tmp330;
  assign tmp332 = decide_ps ? tmp313 : tmp331;
  assign tmp333 = hbusreq1 ? one : zero;
  assign tmp334 = hbusreq0 ? one : zero;
  assign tmp335 = hgrant1_ps ? tmp333 : tmp334;
  assign tmp336 = hmaster0_ps ? tmp333 : tmp334;
  assign tmp337 = hready_ps ? tmp335 : tmp336;
  assign tmp338 = stateG3_1_ps ? tmp68 : one;
  assign tmp339 = stateG3_2_ps ? one : tmp338;
  assign tmp340 = stateA1_ps ? one : tmp339;
  assign tmp341 = hbusreq0 ? tmp340 : one;
  assign tmp342 = stateG3_1_ps ? tmp0 : tmp65;
  assign tmp343 = stateG3_2_ps ? tmp0 : tmp342;
  assign tmp344 = stateG3_1_ps ? tmp2 : tmp68;
  assign tmp345 = stateG3_2_ps ? tmp2 : tmp344;
  assign tmp346 = ~tmp345;
  assign tmp347 = hburst0_ps ? tmp343 : tmp346;
  assign tmp348 = hburst0_ps ? tmp343 : zero;
  assign tmp349 = hburst1_ps ? tmp347 : tmp348;
  assign tmp350 = ~tmp349;
  assign tmp351 = stateA1_ps ? one : tmp350;
  assign tmp352 = hbusreq0 ? tmp351 : one;
  assign tmp353 = hlock1 ? tmp341 : tmp352;
  assign tmp354 = hburst1_ps ? tmp72 : tmp67;
  assign tmp355 = stateG2_ps ? tmp0 : tmp354;
  assign tmp356 = hburst1_ps ? tmp347 : tmp343;
  assign tmp357 = stateA1_ps ? tmp355 : tmp356;
  assign tmp358 = hbusreq0 ? tmp357 : zero;
  assign tmp359 = ~tmp358;
  assign tmp360 = hbusreq1 ? tmp353 : tmp359;
  assign tmp361 = stateA1_ps ? one : tmp1;
  assign tmp362 = ~tmp172;
  assign tmp363 = stateA1_ps ? one : tmp362;
  assign tmp364 = hbusreq0 ? tmp363 : one;
  assign tmp365 = hlock1 ? tmp361 : tmp364;
  assign tmp366 = stateA1_ps ? tmp355 : tmp354;
  assign tmp367 = hbusreq0 ? tmp366 : zero;
  assign tmp368 = ~tmp367;
  assign tmp369 = hbusreq1 ? tmp365 : tmp368;
  assign tmp370 = hready ? tmp360 : tmp369;
  assign tmp371 = locked_ps ? tmp370 : one;
  assign tmp372 = hlock1_ps ? tmp371 : one;
  assign tmp373 = hburst0_ps ? tmp339 : one;
  assign tmp374 = hburst1_ps ? tmp339 : tmp373;
  assign tmp375 = stateA1_ps ? one : tmp374;
  assign tmp376 = hbusreq0 ? tmp375 : one;
  assign tmp377 = hburst0_ps ? tmp339 : tmp295;
  assign tmp378 = hburst1_ps ? tmp339 : tmp377;
  assign tmp379 = ~tmp378;
  assign tmp380 = stateA1_ps ? tmp299 : tmp379;
  assign tmp381 = hbusreq0 ? tmp380 : zero;
  assign tmp382 = ~tmp381;
  assign tmp383 = hbusreq1 ? tmp376 : tmp382;
  assign tmp384 = stateA1_ps ? tmp299 : tmp298;
  assign tmp385 = hbusreq0 ? tmp384 : zero;
  assign tmp386 = ~tmp385;
  assign tmp387 = hbusreq1 ? one : tmp386;
  assign tmp388 = hready ? tmp383 : tmp387;
  assign tmp389 = locked_ps ? tmp388 : one;
  assign tmp390 = hlock1_ps ? tmp389 : one;
  assign tmp391 = hlock0_ps ? tmp372 : tmp390;
  assign tmp392 = hbusreq0_ps ? tmp391 : one;
  assign tmp393 = jx_1_ps ? tmp392 : one;
  assign tmp394 = jx_0_ps ? one : tmp393;
  assign tmp395 = stateA1_ps ? tmp57 : one;
  assign tmp396 = hbusreq0 ? tmp395 : one;
  assign tmp397 = locked_ps ? one : tmp396;
  assign tmp398 = hlock0_ps ? tmp397 : one;
  assign tmp399 = hbusreq0_ps ? tmp398 : one;
  assign tmp400 = jx_1_ps ? tmp399 : one;
  assign tmp401 = jx_0_ps ? one : tmp400;
  assign tmp402 = hbusreq1_ps ? tmp394 : tmp401;
  assign tmp403 = hmaster0_ps ? tmp402 : one;
  assign tmp404 = hburst0_ps ? tmp68 : one;
  assign tmp405 = hburst1_ps ? tmp68 : tmp404;
  assign tmp406 = stateA1_ps ? one : tmp405;
  assign tmp407 = hburst0_ps ? tmp65 : tmp343;
  assign tmp408 = ~tmp407;
  assign tmp409 = hburst1_ps ? tmp68 : tmp408;
  assign tmp410 = ~tmp409;
  assign tmp411 = stateA1_ps ? tmp355 : tmp410;
  assign tmp412 = ~tmp411;
  assign tmp413 = hbusreq0 ? tmp406 : tmp412;
  assign tmp414 = ~tmp357;
  assign tmp415 = hbusreq0 ? tmp351 : tmp414;
  assign tmp416 = hlock1 ? tmp413 : tmp415;
  assign tmp417 = hbusreq1 ? tmp416 : one;
  assign tmp418 = ~tmp366;
  assign tmp419 = hbusreq0 ? tmp363 : tmp418;
  assign tmp420 = hbusreq1 ? tmp419 : one;
  assign tmp421 = hready ? tmp417 : tmp420;
  assign tmp422 = locked_ps ? tmp421 : one;
  assign tmp423 = hburst0_ps ? tmp65 : tmp63;
  assign tmp424 = ~tmp423;
  assign tmp425 = hburst1_ps ? tmp68 : tmp424;
  assign tmp426 = ~tmp425;
  assign tmp427 = stateA1_ps ? tmp299 : tmp426;
  assign tmp428 = ~tmp427;
  assign tmp429 = hbusreq0 ? tmp375 : tmp428;
  assign tmp430 = hbusreq1 ? tmp429 : one;
  assign tmp431 = ~tmp384;
  assign tmp432 = hbusreq0 ? one : tmp431;
  assign tmp433 = hbusreq1 ? tmp432 : one;
  assign tmp434 = hready ? tmp430 : tmp433;
  assign tmp435 = locked_ps ? tmp434 : one;
  assign tmp436 = hlock1_ps ? tmp422 : tmp435;
  assign tmp437 = stateA1_ps ? one : zero;
  assign tmp438 = hbusreq1 ? tmp437 : zero;
  assign tmp439 = ~tmp438;
  assign tmp440 = locked_ps ? one : tmp439;
  assign tmp441 = busreq_ps ? one : tmp440;
  assign tmp442 = hlock1_ps ? tmp441 : one;
  assign tmp443 = hlock0_ps ? tmp436 : tmp442;
  assign tmp444 = jx_1_ps ? tmp443 : one;
  assign tmp445 = jx_0_ps ? tmp444 : one;
  assign tmp446 = hbusreq1_ps ? tmp445 : one;
  assign tmp447 = hmaster0_ps ? one : tmp446;
  assign tmp448 = hgrant1_ps ? tmp403 : tmp447;
  assign tmp449 = stateA1_ps ? one : tmp7;
  assign tmp450 = hbusreq0 ? tmp449 : one;
  assign tmp451 = hlock1 ? tmp450 : tmp364;
  assign tmp452 = hbusreq1 ? tmp451 : tmp368;
  assign tmp453 = stateG3_1_ps ? tmp63 : tmp65;
  assign tmp454 = stateG3_2_ps ? tmp0 : tmp453;
  assign tmp455 = stateG3_1_ps ? one : tmp68;
  assign tmp456 = stateG3_2_ps ? tmp2 : tmp455;
  assign tmp457 = ~tmp456;
  assign tmp458 = hburst0_ps ? tmp454 : tmp457;
  assign tmp459 = hburst0_ps ? tmp454 : zero;
  assign tmp460 = hburst1_ps ? tmp458 : tmp459;
  assign tmp461 = ~tmp460;
  assign tmp462 = stateA1_ps ? one : tmp461;
  assign tmp463 = hbusreq0 ? tmp462 : one;
  assign tmp464 = hlock1 ? tmp361 : tmp463;
  assign tmp465 = hburst1_ps ? tmp458 : tmp454;
  assign tmp466 = stateG2_ps ? tmp0 : tmp465;
  assign tmp467 = stateA1_ps ? tmp466 : tmp465;
  assign tmp468 = hbusreq0 ? tmp467 : zero;
  assign tmp469 = ~tmp468;
  assign tmp470 = hbusreq1 ? tmp464 : tmp469;
  assign tmp471 = hready ? tmp452 : tmp470;
  assign tmp472 = hlock1_ps ? tmp471 : one;
  assign tmp473 = hburst0_ps ? tmp5 : one;
  assign tmp474 = hburst1_ps ? tmp5 : tmp473;
  assign tmp475 = stateA1_ps ? one : tmp474;
  assign tmp476 = hbusreq0 ? tmp475 : one;
  assign tmp477 = stateG3_1_ps ? tmp64 : tmp63;
  assign tmp478 = ~tmp477;
  assign tmp479 = hburst1_ps ? tmp4 : tmp478;
  assign tmp480 = ~tmp479;
  assign tmp481 = stateG2_ps ? tmp0 : tmp480;
  assign tmp482 = stateG3_2_ps ? tmp63 : tmp477;
  assign tmp483 = ~tmp482;
  assign tmp484 = hburst0_ps ? tmp5 : tmp483;
  assign tmp485 = hburst1_ps ? tmp5 : tmp484;
  assign tmp486 = ~tmp485;
  assign tmp487 = stateA1_ps ? tmp481 : tmp486;
  assign tmp488 = hbusreq0 ? tmp487 : zero;
  assign tmp489 = ~tmp488;
  assign tmp490 = hbusreq1 ? tmp476 : tmp489;
  assign tmp491 = hready ? tmp490 : tmp387;
  assign tmp492 = hlock1_ps ? tmp491 : one;
  assign tmp493 = hlock0_ps ? tmp472 : tmp492;
  assign tmp494 = hbusreq0_ps ? tmp493 : one;
  assign tmp495 = jx_1_ps ? tmp494 : one;
  assign tmp496 = jx_0_ps ? one : tmp495;
  assign tmp497 = hbusreq1_ps ? tmp496 : one;
  assign tmp498 = hburst0_ps ? tmp4 : one;
  assign tmp499 = hburst1_ps ? tmp4 : tmp498;
  assign tmp500 = stateA1_ps ? one : tmp499;
  assign tmp501 = hburst0_ps ? tmp477 : tmp67;
  assign tmp502 = ~tmp501;
  assign tmp503 = hburst1_ps ? tmp4 : tmp502;
  assign tmp504 = ~tmp503;
  assign tmp505 = stateA1_ps ? tmp355 : tmp504;
  assign tmp506 = ~tmp505;
  assign tmp507 = hbusreq0 ? tmp500 : tmp506;
  assign tmp508 = hlock1 ? tmp507 : tmp419;
  assign tmp509 = hbusreq1 ? tmp508 : one;
  assign tmp510 = ~tmp467;
  assign tmp511 = hbusreq0 ? tmp462 : tmp510;
  assign tmp512 = hbusreq1 ? tmp511 : one;
  assign tmp513 = hready ? tmp509 : tmp512;
  assign tmp514 = stateA1_ps ? tmp481 : tmp480;
  assign tmp515 = ~tmp514;
  assign tmp516 = hbusreq0 ? tmp475 : tmp515;
  assign tmp517 = hbusreq1 ? tmp516 : one;
  assign tmp518 = hready ? tmp517 : tmp433;
  assign tmp519 = hlock1_ps ? tmp513 : tmp518;
  assign tmp520 = hlock0_ps ? tmp519 : one;
  assign tmp521 = jx_1_ps ? tmp520 : one;
  assign tmp522 = jx_0_ps ? tmp521 : one;
  assign tmp523 = hbusreq1_ps ? tmp522 : one;
  assign tmp524 = hmaster0_ps ? tmp497 : tmp523;
  assign tmp525 = hready_ps ? tmp448 : tmp524;
  assign tmp526 = ~tmp344;
  assign tmp527 = hburst0_ps ? tmp342 : tmp526;
  assign tmp528 = hburst0_ps ? tmp342 : zero;
  assign tmp529 = hburst1_ps ? tmp527 : tmp528;
  assign tmp530 = ~tmp529;
  assign tmp531 = stateA1_ps ? one : tmp530;
  assign tmp532 = hbusreq0 ? tmp531 : one;
  assign tmp533 = hburst0_ps ? tmp342 : tmp343;
  assign tmp534 = hburst1_ps ? tmp527 : tmp533;
  assign tmp535 = stateA1_ps ? tmp355 : tmp534;
  assign tmp536 = hbusreq0 ? tmp535 : zero;
  assign tmp537 = ~tmp536;
  assign tmp538 = hbusreq1 ? tmp532 : tmp537;
  assign tmp539 = hburst0_ps ? tmp63 : tmp67;
  assign tmp540 = ~tmp539;
  assign tmp541 = hburst1_ps ? one : tmp540;
  assign tmp542 = ~tmp541;
  assign tmp543 = stateA1_ps ? tmp355 : tmp542;
  assign tmp544 = hbusreq0 ? tmp543 : zero;
  assign tmp545 = ~tmp544;
  assign tmp546 = hbusreq1 ? one : tmp545;
  assign tmp547 = hready ? tmp538 : tmp546;
  assign tmp548 = hbusreq1 ? tmp59 : zero;
  assign tmp549 = ~tmp361;
  assign tmp550 = hbusreq1 ? tmp114 : tmp549;
  assign tmp551 = hready ? tmp548 : tmp550;
  assign tmp552 = locked_ps ? tmp547 : tmp551;
  assign tmp553 = ~tmp69;
  assign tmp554 = hburst0_ps ? tmp66 : tmp553;
  assign tmp555 = stateG2_ps ? tmp0 : tmp554;
  assign tmp556 = stateA1_ps ? tmp555 : tmp529;
  assign tmp557 = hbusreq0 ? tmp556 : zero;
  assign tmp558 = stateA1_ps ? tmp555 : tmp534;
  assign tmp559 = hbusreq0 ? tmp558 : zero;
  assign tmp560 = hbusreq1 ? tmp557 : tmp559;
  assign tmp561 = stateA1_ps ? tmp555 : zero;
  assign tmp562 = hbusreq0 ? tmp561 : zero;
  assign tmp563 = stateA1_ps ? tmp555 : tmp542;
  assign tmp564 = hbusreq0 ? tmp563 : zero;
  assign tmp565 = hbusreq1 ? tmp562 : tmp564;
  assign tmp566 = hready ? tmp560 : tmp565;
  assign tmp567 = stateA1_ps ? one : tmp57;
  assign tmp568 = hbusreq1 ? tmp567 : one;
  assign tmp569 = hready ? tmp568 : tmp361;
  assign tmp570 = locked_ps ? tmp566 : tmp569;
  assign tmp571 = ~tmp570;
  assign tmp572 = busreq_ps ? tmp552 : tmp571;
  assign tmp573 = hbusreq0_ps ? tmp572 : one;
  assign tmp574 = jx_1_ps ? tmp573 : one;
  assign tmp575 = jx_0_ps ? one : tmp574;
  assign tmp576 = hmaster0_ps ? tmp575 : one;
  assign tmp577 = hbusreq1 ? tmp415 : one;
  assign tmp578 = ~tmp543;
  assign tmp579 = hbusreq0 ? one : tmp578;
  assign tmp580 = hbusreq1 ? tmp579 : one;
  assign tmp581 = hready ? tmp577 : tmp580;
  assign tmp582 = hbusreq1 ? tmp59 : tmp114;
  assign tmp583 = hready ? tmp582 : tmp114;
  assign tmp584 = locked_ps ? tmp581 : tmp583;
  assign tmp585 = stateG2_ps ? tmp0 : tmp72;
  assign tmp586 = stateA1_ps ? tmp585 : tmp349;
  assign tmp587 = stateA1_ps ? tmp585 : tmp356;
  assign tmp588 = hbusreq0 ? tmp586 : tmp587;
  assign tmp589 = hbusreq1 ? tmp588 : zero;
  assign tmp590 = stateA1_ps ? tmp585 : zero;
  assign tmp591 = stateA1_ps ? tmp585 : tmp542;
  assign tmp592 = hbusreq0 ? tmp590 : tmp591;
  assign tmp593 = hbusreq1 ? tmp592 : zero;
  assign tmp594 = hready ? tmp589 : tmp593;
  assign tmp595 = hbusreq1 ? tmp567 : tmp115;
  assign tmp596 = hbusreq1 ? tmp361 : tmp115;
  assign tmp597 = hready ? tmp595 : tmp596;
  assign tmp598 = locked_ps ? tmp594 : tmp597;
  assign tmp599 = ~tmp598;
  assign tmp600 = busreq_ps ? tmp584 : tmp599;
  assign tmp601 = jx_1_ps ? tmp600 : one;
  assign tmp602 = jx_0_ps ? tmp601 : one;
  assign tmp603 = hbusreq1_ps ? tmp602 : one;
  assign tmp604 = hmaster0_ps ? one : tmp603;
  assign tmp605 = hgrant1_ps ? tmp576 : tmp604;
  assign tmp606 = hbusreq1 ? tmp364 : tmp368;
  assign tmp607 = stateA1_ps ? tmp0 : one;
  assign tmp608 = hburst1_ps ? tmp122 : tmp118;
  assign tmp609 = stateG2_ps ? one : tmp608;
  assign tmp610 = hburst0_ps ? tmp63 : tmp454;
  assign tmp611 = ~tmp610;
  assign tmp612 = hburst1_ps ? one : tmp611;
  assign tmp613 = ~tmp612;
  assign tmp614 = stateA1_ps ? tmp609 : tmp613;
  assign tmp615 = ~tmp607;
  assign tmp616 = hbusreq0 ? tmp614 : tmp615;
  assign tmp617 = ~tmp616;
  assign tmp618 = hbusreq1 ? tmp607 : tmp617;
  assign tmp619 = hready ? tmp606 : tmp618;
  assign tmp620 = hbusreq1 ? tmp114 : tmp0;
  assign tmp621 = locked_ps ? tmp619 : tmp620;
  assign tmp622 = stateA1_ps ? tmp555 : tmp172;
  assign tmp623 = hbusreq0 ? tmp622 : zero;
  assign tmp624 = stateA1_ps ? tmp555 : tmp354;
  assign tmp625 = hbusreq0 ? tmp624 : zero;
  assign tmp626 = hbusreq1 ? tmp623 : tmp625;
  assign tmp627 = ~tmp119;
  assign tmp628 = hburst0_ps ? tmp117 : tmp627;
  assign tmp629 = stateG2_ps ? one : tmp628;
  assign tmp630 = stateA1_ps ? tmp629 : zero;
  assign tmp631 = hbusreq0 ? tmp630 : tmp615;
  assign tmp632 = stateA1_ps ? tmp629 : tmp613;
  assign tmp633 = hbusreq0 ? tmp632 : tmp615;
  assign tmp634 = hbusreq1 ? tmp631 : tmp633;
  assign tmp635 = hready ? tmp626 : tmp634;
  assign tmp636 = locked_ps ? tmp635 : tmp1;
  assign tmp637 = ~tmp636;
  assign tmp638 = busreq_ps ? tmp621 : tmp637;
  assign tmp639 = hbusreq0_ps ? tmp638 : one;
  assign tmp640 = jx_1_ps ? tmp639 : one;
  assign tmp641 = jx_0_ps ? one : tmp640;
  assign tmp642 = hmaster0_ps ? tmp641 : one;
  assign tmp643 = ~tmp614;
  assign tmp644 = hbusreq0 ? tmp607 : tmp643;
  assign tmp645 = hbusreq1 ? tmp644 : tmp607;
  assign tmp646 = hready ? tmp420 : tmp645;
  assign tmp647 = locked_ps ? tmp646 : tmp114;
  assign tmp648 = stateA1_ps ? tmp585 : tmp172;
  assign tmp649 = stateA1_ps ? tmp585 : tmp354;
  assign tmp650 = hbusreq0 ? tmp648 : tmp649;
  assign tmp651 = hbusreq1 ? tmp650 : zero;
  assign tmp652 = stateG2_ps ? one : tmp122;
  assign tmp653 = stateA1_ps ? tmp652 : zero;
  assign tmp654 = stateA1_ps ? tmp652 : tmp613;
  assign tmp655 = hbusreq0 ? tmp653 : tmp654;
  assign tmp656 = hbusreq1 ? tmp655 : tmp615;
  assign tmp657 = hready ? tmp651 : tmp656;
  assign tmp658 = hbusreq1 ? tmp0 : tmp114;
  assign tmp659 = ~tmp658;
  assign tmp660 = locked_ps ? tmp657 : tmp659;
  assign tmp661 = ~tmp660;
  assign tmp662 = busreq_ps ? tmp647 : tmp661;
  assign tmp663 = jx_1_ps ? tmp662 : one;
  assign tmp664 = jx_0_ps ? tmp663 : one;
  assign tmp665 = hbusreq1_ps ? tmp664 : one;
  assign tmp666 = hmaster0_ps ? one : tmp665;
  assign tmp667 = hgrant1_ps ? tmp642 : tmp666;
  assign tmp668 = hready_ps ? tmp605 : tmp667;
  assign tmp669 = decide_ps ? tmp525 : tmp668;
  assign tmp670 = ~tmp669;
  assign tmp671 = hready_ps ? tmp53 : tmp0;
  assign tmp672 = stateG3_1_ps ? tmp68 : tmp3;
  assign tmp673 = stateG3_2_ps ? one : tmp672;
  assign tmp674 = stateG3_1_ps ? tmp65 : tmp64;
  assign tmp675 = stateG3_2_ps ? tmp63 : tmp674;
  assign tmp676 = ~tmp675;
  assign tmp677 = hburst0_ps ? tmp673 : tmp676;
  assign tmp678 = hburst1_ps ? tmp677 : tmp673;
  assign tmp679 = stateG2_ps ? one : tmp678;
  assign tmp680 = stateG3_1_ps ? tmp2 : one;
  assign tmp681 = stateG3_2_ps ? one : tmp680;
  assign tmp682 = stateG2_ps ? one : tmp681;
  assign tmp683 = hready_ps ? tmp679 : tmp682;
  assign tmp684 = stateA1_ps ? tmp678 : tmp679;
  assign tmp685 = busreq_ps ? tmp679 : tmp684;
  assign tmp686 = jx_1_ps ? tmp679 : tmp685;
  assign tmp687 = jx_0_ps ? tmp679 : tmp686;
  assign tmp688 = stateA1_ps ? tmp681 : tmp682;
  assign tmp689 = busreq_ps ? tmp682 : tmp688;
  assign tmp690 = jx_1_ps ? tmp682 : tmp689;
  assign tmp691 = jx_0_ps ? tmp682 : tmp690;
  assign tmp692 = hready_ps ? tmp687 : tmp691;
  assign tmp693 = decide_ps ? tmp683 : tmp692;
  assign tmp694 = ~tmp693;
  assign tmp695 = stateG2_ps ? one : tmp339;
  assign tmp696 = stateG3_2_ps ? tmp63 : tmp64;
  assign tmp697 = ~tmp696;
  assign tmp698 = hburst0_ps ? tmp7 : tmp697;
  assign tmp699 = hburst1_ps ? tmp698 : tmp7;
  assign tmp700 = stateG2_ps ? one : tmp699;
  assign tmp701 = hready_ps ? tmp695 : tmp700;
  assign tmp702 = stateA1_ps ? tmp339 : tmp695;
  assign tmp703 = busreq_ps ? tmp695 : tmp702;
  assign tmp704 = jx_1_ps ? tmp695 : tmp703;
  assign tmp705 = jx_0_ps ? tmp695 : tmp704;
  assign tmp706 = stateA1_ps ? tmp699 : tmp700;
  assign tmp707 = busreq_ps ? tmp700 : tmp706;
  assign tmp708 = jx_1_ps ? tmp700 : tmp707;
  assign tmp709 = jx_0_ps ? tmp700 : tmp708;
  assign tmp710 = hready_ps ? tmp705 : tmp709;
  assign tmp711 = decide_ps ? tmp701 : tmp710;
  assign tmp712 = ~tmp711;
  assign tmp713 = hburst0_ps ? one : tmp1;
  assign tmp714 = hburst1_ps ? one : tmp713;
  assign tmp715 = ~tmp714;
  assign tmp716 = stateA1_ps ? one : tmp715;
  assign tmp717 = ~tmp567;
  assign tmp718 = hbusreq1_ps ? tmp716 : tmp717;
  assign tmp719 = busreq_ps ? tmp59 : tmp717;
  assign tmp720 = hlock0_ps ? tmp59 : tmp719;
  assign tmp721 = jx_1_ps ? tmp719 : tmp720;
  assign tmp722 = hbusreq0_ps ? tmp59 : tmp717;
  assign tmp723 = jx_0_ps ? tmp721 : tmp722;
  assign tmp724 = hbusreq1_ps ? tmp723 : tmp722;
  assign tmp725 = hmaster0_ps ? tmp718 : tmp724;
  assign tmp726 = hlock0_ps ? one : tmp567;
  assign tmp727 = hbusreq0_ps ? tmp726 : tmp567;
  assign tmp728 = jx_1_ps ? tmp727 : tmp726;
  assign tmp729 = jx_0_ps ? tmp726 : tmp728;
  assign tmp730 = ~tmp729;
  assign tmp731 = hbusreq1_ps ? tmp59 : tmp730;
  assign tmp732 = hlock0_ps ? tmp716 : tmp719;
  assign tmp733 = hlock0_ps ? tmp716 : tmp59;
  assign tmp734 = hbusreq0_ps ? tmp733 : tmp717;
  assign tmp735 = jx_1_ps ? tmp734 : tmp732;
  assign tmp736 = jx_0_ps ? tmp732 : tmp735;
  assign tmp737 = stateA1_ps ? tmp0 : tmp715;
  assign tmp738 = hlock0_ps ? tmp737 : tmp719;
  assign tmp739 = hlock0_ps ? tmp737 : tmp59;
  assign tmp740 = hbusreq0_ps ? tmp739 : tmp717;
  assign tmp741 = jx_1_ps ? tmp740 : tmp738;
  assign tmp742 = jx_0_ps ? tmp738 : tmp741;
  assign tmp743 = hbusreq1_ps ? tmp736 : tmp742;
  assign tmp744 = hmaster0_ps ? tmp731 : tmp743;
  assign tmp745 = hgrant1_ps ? tmp725 : tmp744;
  assign tmp746 = jx_0_ps ? tmp732 : tmp734;
  assign tmp747 = hbusreq1_ps ? tmp746 : tmp734;
  assign tmp748 = hmaster0_ps ? tmp718 : tmp747;
  assign tmp749 = ~tmp727;
  assign tmp750 = hbusreq1_ps ? tmp716 : tmp749;
  assign tmp751 = hbusreq1_ps ? tmp746 : tmp740;
  assign tmp752 = hmaster0_ps ? tmp750 : tmp751;
  assign tmp753 = hgrant1_ps ? tmp748 : tmp752;
  assign tmp754 = hready_ps ? tmp745 : tmp753;
  assign tmp755 = stateA1_ps ? one : tmp714;
  assign tmp756 = ~tmp755;
  assign tmp757 = busreq_ps ? tmp716 : tmp756;
  assign tmp758 = jx_1_ps ? tmp716 : tmp757;
  assign tmp759 = jx_0_ps ? tmp758 : tmp757;
  assign tmp760 = ~tmp757;
  assign tmp761 = jx_1_ps ? tmp755 : tmp760;
  assign tmp762 = jx_0_ps ? tmp761 : tmp760;
  assign tmp763 = ~tmp762;
  assign tmp764 = hbusreq1_ps ? tmp759 : tmp763;
  assign tmp765 = jx_1_ps ? tmp722 : tmp719;
  assign tmp766 = jx_0_ps ? tmp719 : tmp765;
  assign tmp767 = hmaster0_ps ? tmp764 : tmp766;
  assign tmp768 = hbusreq1_ps ? tmp59 : tmp717;
  assign tmp769 = hbusreq0_ps ? tmp716 : tmp756;
  assign tmp770 = jx_1_ps ? tmp769 : tmp757;
  assign tmp771 = jx_0_ps ? tmp757 : tmp770;
  assign tmp772 = hmaster0_ps ? tmp768 : tmp771;
  assign tmp773 = hgrant1_ps ? tmp767 : tmp772;
  assign tmp774 = decide_ps ? tmp754 : tmp773;
  assign tmp775 = hbusreq1_ps ? one : zero;
  assign tmp776 = hgrant1_ps ? one : tmp775;
  assign tmp777 = ~tmp776;
  assign tmp778 = jx_1_ps ? tmp185 : tmp437;
  assign tmp779 = jx_0_ps ? tmp274 : tmp778;
  assign tmp780 = ~tmp437;
  assign tmp781 = jx_1_ps ? one : tmp780;
  assign tmp782 = jx_0_ps ? tmp256 : tmp781;
  assign tmp783 = ~tmp781;
  assign tmp784 = jx_0_ps ? tmp274 : tmp783;
  assign tmp785 = ~tmp784;
  assign tmp786 = hbusreq1_ps ? tmp782 : tmp785;
  assign tmp787 = ~tmp786;
  assign tmp788 = hmaster0_ps ? tmp779 : tmp787;
  assign tmp789 = ~tmp788;
  assign hmaster0 = tmp160;
  assign hmastlock = tmp671;
  assign start = tmp168;
  assign decide = tmp670;
  assign locked = tmp157;
  assign hgrant0 = tmp252;
  assign hgrant1 = tmp241;
  assign busreq = tmp337;
  assign stateA1 = tmp774;
  assign stateG2 = tmp332;
  assign stateG2_0 = zero;
  assign stateG2_1 = zero;
  assign stateG3_0 = tmp712;
  assign stateG3_1 = tmp694;
  assign stateG3_2 = tmp51;
  assign stateG10_1 = tmp777;
  assign jx_0 = tmp789;
  assign jx_1 = tmp294;
  assign zero = 0;
  assign one = 1;
  initial
  begin
    hready_ps = 0;
    hbusreq0_ps = 0;
    hlock0_ps = 0;
    hbusreq1_ps = 0;
    hlock1_ps = 0;
    hburst0_ps = 0;
    hburst1_ps = 0;
    hmaster0_ps = 0;
    hmastlock_ps = 0;
    start_ps = 1;
    decide_ps = 1;
    locked_ps = 0;
    hgrant0_ps = 1;
    hgrant1_ps = 0;
    busreq_ps = 0;
    stateA1_ps = 0;
    stateG2_ps = 0;
    stateG2_0_ps = 0;
    stateG2_1_ps = 0;
    stateG3_0_ps = 0;
    stateG3_1_ps = 0;
    stateG3_2_ps = 0;
    stateG10_1_ps = 0;
    jx_0_ps = 0;
    jx_1_ps = 0;
  end
  always @(posedge clock)
  begin
    hready_ps = hready;
    hbusreq0_ps = hbusreq0;
    hlock0_ps = hlock0;
    hbusreq1_ps = hbusreq1;
    hlock1_ps = hlock1;
    hburst0_ps = hburst0;
    hburst1_ps = hburst1;
    hmaster0_ps = tmp160;
    hmastlock_ps = tmp671;
    start_ps = tmp168;
    decide_ps = tmp670;
    locked_ps = tmp157;
    hgrant0_ps = tmp252;
    hgrant1_ps = tmp241;
    busreq_ps = tmp337;
    stateA1_ps = tmp774;
    stateG2_ps = tmp332;
    stateG2_0_ps = zero;
    stateG2_1_ps = zero;
    stateG3_0_ps = tmp712;
    stateG3_1_ps = tmp694;
    stateG3_2_ps = tmp51;
    stateG10_1_ps = tmp777;
    jx_0_ps = tmp789;
    jx_1_ps = tmp294;
  end
endmodule

